package monitor_piso;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	import sequence_item_piso::*;

	class monitor_piso extends uvm_monitor;
		`uvm_component_utils(monitor_piso)

		virtual piso_if  vif;
		uvm_analysis_port #(sequence_item_piso) item_collected_port;

		function new(string name, uvm_component parent);
			super.new(name, parent);
		endfunction : new

        function void connect_phase(uvm_phase phase);
            if (!uvm_config_db#(virtual piso_if)::get(this,"","piso_if", vif))
	            `uvm_error("NOVIF",{"virtual interface must be set for: ",get_full_name(),".vif"})
		endfunction: connect_phase

		virtual function void build_phase(uvm_phase phase);
			super.build_phase(phase);
			item_collected_port = new("item_collected_port", this);
		endfunction : build_phase

		virtual task run_phase(uvm_phase phase);
			super.run_phase(phase);
			forever begin
				sample_item();
			end
		endtask : run_phase

		virtual task sample_item();
			sequence_item_piso resp = sequence_item_piso::type_id::create("resp");            
			@(posedge vif.BitCLK);
            //***************************//
            // TODO: Sample Outputs Here //
			logic [9:0] expected_data;
        logic [9:0] temp_reg;
        int i;

        // Process serial data and compare with expected output
        forever begin
            @(posedge vif.BitCLK);
            if (vif.Reset == 0) begin
                // Reset: expected data should be 0
                expected_data = 10'b0;
                temp_reg = 10'b0;
            end else begin
                // Shift expected data by one position
                expected_data = expected_data >> 1;
                expected_data[9] = vif.TxParallel_10[9]; // shift in the first bit of parallel data
                temp_reg = expected_data;
                ap_serial.write(vif.Serial); // Send serial output for analysis
            end
            //***************************//
			// example: resp.signal = vif.signal
			item_collected_port.write(resp);
		end
		endtask : sample_item

	endclass 
endpackage