module assertions_cdr_top (cdr_top_if.DUT _if);
    
    //*****************************//
    // TODO: Write Assertions Here //
    //*****************************//

endmodule