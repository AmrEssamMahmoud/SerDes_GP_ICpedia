module assertions_equalization_top (equalization_top_if.DUT _if);
    
    //*****************************//
    // TODO: Write Assertions Here //
    //*****************************//

endmodule