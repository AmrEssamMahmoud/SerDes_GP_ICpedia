module assertions_buffer (buffer_if.DUT _if);
    
    // assertion for wrtite and read pointer incrementation 
    // assertion for read and write pointer for stalltion in case of skp and for installtion in case of read while empty and write while full
    // assertion for full and empty flags
    // assertion for reset

    //*****************************//
    // TODO: Write Assertions Here //
    //*****************************//

endmodule