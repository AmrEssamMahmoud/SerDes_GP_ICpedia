module channel (
    input in,
    output out
);

    assign out = in;

endmodule