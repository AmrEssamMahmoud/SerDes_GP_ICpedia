module equalizer (
    input in,
    output out
);

    assign out = in;

endmodule